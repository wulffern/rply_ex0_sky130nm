magic
tech sky130B
magscale 1 2
timestamp 1671570105
<< locali >>
rect 3260 740 3360 1120
rect 3640 740 3740 1120
rect 3960 740 4060 1120
rect 4340 740 4440 1120
rect 4660 740 4760 1120
rect 5040 740 5140 1120
rect 5360 740 5460 1120
rect 5740 740 5840 1120
rect 6060 740 6160 1120
rect 6440 740 6540 1120
rect 6760 740 6860 1120
rect 7140 740 7240 1120
rect 3280 400 3720 440
rect 3980 400 4420 440
rect 4680 400 5120 440
rect 5380 400 5820 440
rect 6080 400 6520 440
rect 6800 400 7240 440
rect 3200 300 7300 400
<< metal1 >>
rect 3400 1360 7290 1420
rect 4870 1300 4930 1360
rect 3460 1060 3540 1300
rect 4160 1060 4240 1300
rect 4154 980 4160 1060
rect 4240 980 4246 1060
rect 3460 640 3540 980
rect 4160 640 4240 980
rect 4860 640 4940 1300
rect 5560 1060 5640 1300
rect 6260 1060 6340 1300
rect 5554 980 5560 1060
rect 5640 980 5646 1060
rect 5560 640 5640 980
rect 6260 640 6340 980
rect 6960 1060 7040 1300
rect 6960 640 7040 980
rect 3400 520 7290 580
<< via1 >>
rect 3460 980 3540 1060
rect 4160 980 4240 1060
rect 5560 980 5640 1060
rect 6260 980 6340 1060
rect 6960 980 7040 1060
<< metal2 >>
rect 4160 1060 4240 1066
rect 5560 1060 5640 1066
rect 3454 980 3460 1060
rect 3540 980 4160 1060
rect 4240 980 5560 1060
rect 5640 980 6260 1060
rect 6340 980 6960 1060
rect 7040 980 7220 1060
rect 4160 974 4240 980
rect 5560 974 5640 980
use sky130_fd_pr__nfet_01v8_5CE34N  sky130_fd_pr__nfet_01v8_5CE34N_0
timestamp 1671548393
transform 1 0 6997 0 1 970
box -297 -570 297 570
use sky130_fd_pr__nfet_01v8_5CE34N  sky130_fd_pr__nfet_01v8_5CE34N_1
timestamp 1671548393
transform 1 0 3497 0 1 970
box -297 -570 297 570
use sky130_fd_pr__nfet_01v8_5CE34N  sky130_fd_pr__nfet_01v8_5CE34N_2
timestamp 1671548393
transform 1 0 4197 0 1 970
box -297 -570 297 570
use sky130_fd_pr__nfet_01v8_5CE34N  sky130_fd_pr__nfet_01v8_5CE34N_3
timestamp 1671548393
transform 1 0 4897 0 1 970
box -297 -570 297 570
use sky130_fd_pr__nfet_01v8_5CE34N  sky130_fd_pr__nfet_01v8_5CE34N_4
timestamp 1671548393
transform 1 0 5597 0 1 970
box -297 -570 297 570
use sky130_fd_pr__nfet_01v8_5CE34N  sky130_fd_pr__nfet_01v8_5CE34N_5
timestamp 1671548393
transform 1 0 6297 0 1 970
box -297 -570 297 570
<< labels >>
flabel metal1 4460 1360 4520 1420 0 FreeSans 320 0 0 0 IBPS_4U
port 2 nsew
flabel locali 4200 300 4280 380 0 FreeSans 320 0 0 0 VSS
port 1 nsew
flabel metal2 4520 980 4600 1060 0 FreeSans 320 0 0 0 IBNS_20U
port 3 nsew
<< end >>
